module stage_execute();
endmodule