module stage_memory();
endmodule