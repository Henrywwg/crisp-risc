module memory(
    input clk,
    input rst_n,
    input 
);



endmodule