module stage_writeback();
endmodule