module reg_file(clk, rst_n, );


endmodule